** Profile: "SCHEMATIC1-monofasicoduplicadordetension1"  [ C:\Users\emile\Desktop\practica 1 ,1-PSpiceFiles\3\monofasico duplicador de tension-PSpiceFiles\SCHEMATIC1\monofasicoduplicadordetension1.sim ] 

** Creating circuit file "monofasicoduplicadordetension1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 100m 40m 100m 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
