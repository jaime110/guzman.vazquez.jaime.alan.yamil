** Profile: "SCHEMATIC1-TENSIONDESALIDA"  [ C:\Users\emile\Desktop\practica 1 ,1-PSpiceFiles\6\monofasico duplicador de tension-PSpiceFiles\SCHEMATIC1\TENSIONDESALIDA.sim ] 

** Creating circuit file "TENSIONDESALIDA.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 40m 0 40m 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
